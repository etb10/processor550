module lab(
	input[4:0] register_index,
	input[31:0] threshold_value,
	input[31:0] incrementer_value,
	input initialize_WE,
	input increase_address,
	input clock,
	input reset,
	output[31:0] address_out,
	output loop
	);



endmodule // lab